
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_LINEAR.weights_stream_V_V_0_U.if_read;
    assign fifo_intf_1.wr_en = AESL_inst_LINEAR.weights_stream_V_V_0_U.if_write;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_0_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0_blk_n);
    assign fifo_intf_1.finish = finish;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_LINEAR.weights_stream_V_V_1_U.if_read;
    assign fifo_intf_2.wr_en = AESL_inst_LINEAR.weights_stream_V_V_1_U.if_write;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_01_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_071_blk_n);
    assign fifo_intf_2.finish = finish;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_LINEAR.weights_stream_V_V_2_U.if_read;
    assign fifo_intf_3.wr_en = AESL_inst_LINEAR.weights_stream_V_V_2_U.if_write;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_02_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_072_blk_n);
    assign fifo_intf_3.finish = finish;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_LINEAR.weights_stream_V_V_3_U.if_read;
    assign fifo_intf_4.wr_en = AESL_inst_LINEAR.weights_stream_V_V_3_U.if_write;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_03_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_073_blk_n);
    assign fifo_intf_4.finish = finish;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_LINEAR.weights_stream_V_V_4_U.if_read;
    assign fifo_intf_5.wr_en = AESL_inst_LINEAR.weights_stream_V_V_4_U.if_write;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_04_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_074_blk_n);
    assign fifo_intf_5.finish = finish;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_LINEAR.weights_stream_V_V_5_U.if_read;
    assign fifo_intf_6.wr_en = AESL_inst_LINEAR.weights_stream_V_V_5_U.if_write;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_05_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_075_blk_n);
    assign fifo_intf_6.finish = finish;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_LINEAR.weights_stream_V_V_6_U.if_read;
    assign fifo_intf_7.wr_en = AESL_inst_LINEAR.weights_stream_V_V_6_U.if_write;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_06_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_076_blk_n);
    assign fifo_intf_7.finish = finish;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_LINEAR.weights_stream_V_V_7_U.if_read;
    assign fifo_intf_8.wr_en = AESL_inst_LINEAR.weights_stream_V_V_7_U.if_write;
    assign fifo_intf_8.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_07_blk_n);
    assign fifo_intf_8.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_077_blk_n);
    assign fifo_intf_8.finish = finish;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_LINEAR.weights_stream_V_V_8_U.if_read;
    assign fifo_intf_9.wr_en = AESL_inst_LINEAR.weights_stream_V_V_8_U.if_write;
    assign fifo_intf_9.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_08_blk_n);
    assign fifo_intf_9.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_078_blk_n);
    assign fifo_intf_9.finish = finish;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_LINEAR.weights_stream_V_V_9_U.if_read;
    assign fifo_intf_10.wr_en = AESL_inst_LINEAR.weights_stream_V_V_9_U.if_write;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_09_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_079_blk_n);
    assign fifo_intf_10.finish = finish;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_LINEAR.weights_stream_V_V_10_U.if_read;
    assign fifo_intf_11.wr_en = AESL_inst_LINEAR.weights_stream_V_V_10_U.if_write;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_010_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_080_blk_n);
    assign fifo_intf_11.finish = finish;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_LINEAR.weights_stream_V_V_11_U.if_read;
    assign fifo_intf_12.wr_en = AESL_inst_LINEAR.weights_stream_V_V_11_U.if_write;
    assign fifo_intf_12.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_011_blk_n);
    assign fifo_intf_12.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_081_blk_n);
    assign fifo_intf_12.finish = finish;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_LINEAR.weights_stream_V_V_12_U.if_read;
    assign fifo_intf_13.wr_en = AESL_inst_LINEAR.weights_stream_V_V_12_U.if_write;
    assign fifo_intf_13.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_012_blk_n);
    assign fifo_intf_13.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_082_blk_n);
    assign fifo_intf_13.finish = finish;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_LINEAR.weights_stream_V_V_13_U.if_read;
    assign fifo_intf_14.wr_en = AESL_inst_LINEAR.weights_stream_V_V_13_U.if_write;
    assign fifo_intf_14.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_013_blk_n);
    assign fifo_intf_14.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_083_blk_n);
    assign fifo_intf_14.finish = finish;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_LINEAR.weights_stream_V_V_14_U.if_read;
    assign fifo_intf_15.wr_en = AESL_inst_LINEAR.weights_stream_V_V_14_U.if_write;
    assign fifo_intf_15.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_014_blk_n);
    assign fifo_intf_15.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_084_blk_n);
    assign fifo_intf_15.finish = finish;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_LINEAR.weights_stream_V_V_15_U.if_read;
    assign fifo_intf_16.wr_en = AESL_inst_LINEAR.weights_stream_V_V_15_U.if_write;
    assign fifo_intf_16.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_015_blk_n);
    assign fifo_intf_16.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_085_blk_n);
    assign fifo_intf_16.finish = finish;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_LINEAR.weights_stream_V_V_16_U.if_read;
    assign fifo_intf_17.wr_en = AESL_inst_LINEAR.weights_stream_V_V_16_U.if_write;
    assign fifo_intf_17.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_016_blk_n);
    assign fifo_intf_17.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_086_blk_n);
    assign fifo_intf_17.finish = finish;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_LINEAR.weights_stream_V_V_17_U.if_read;
    assign fifo_intf_18.wr_en = AESL_inst_LINEAR.weights_stream_V_V_17_U.if_write;
    assign fifo_intf_18.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_017_blk_n);
    assign fifo_intf_18.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_087_blk_n);
    assign fifo_intf_18.finish = finish;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_LINEAR.weights_stream_V_V_18_U.if_read;
    assign fifo_intf_19.wr_en = AESL_inst_LINEAR.weights_stream_V_V_18_U.if_write;
    assign fifo_intf_19.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_018_blk_n);
    assign fifo_intf_19.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_088_blk_n);
    assign fifo_intf_19.finish = finish;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_LINEAR.weights_stream_V_V_19_U.if_read;
    assign fifo_intf_20.wr_en = AESL_inst_LINEAR.weights_stream_V_V_19_U.if_write;
    assign fifo_intf_20.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_019_blk_n);
    assign fifo_intf_20.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_089_blk_n);
    assign fifo_intf_20.finish = finish;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_LINEAR.weights_stream_V_V_20_U.if_read;
    assign fifo_intf_21.wr_en = AESL_inst_LINEAR.weights_stream_V_V_20_U.if_write;
    assign fifo_intf_21.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_020_blk_n);
    assign fifo_intf_21.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_090_blk_n);
    assign fifo_intf_21.finish = finish;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_LINEAR.weights_stream_V_V_21_U.if_read;
    assign fifo_intf_22.wr_en = AESL_inst_LINEAR.weights_stream_V_V_21_U.if_write;
    assign fifo_intf_22.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_021_blk_n);
    assign fifo_intf_22.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_091_blk_n);
    assign fifo_intf_22.finish = finish;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_LINEAR.weights_stream_V_V_22_U.if_read;
    assign fifo_intf_23.wr_en = AESL_inst_LINEAR.weights_stream_V_V_22_U.if_write;
    assign fifo_intf_23.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_022_blk_n);
    assign fifo_intf_23.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_092_blk_n);
    assign fifo_intf_23.finish = finish;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_LINEAR.weights_stream_V_V_23_U.if_read;
    assign fifo_intf_24.wr_en = AESL_inst_LINEAR.weights_stream_V_V_23_U.if_write;
    assign fifo_intf_24.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_023_blk_n);
    assign fifo_intf_24.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_093_blk_n);
    assign fifo_intf_24.finish = finish;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_LINEAR.weights_stream_V_V_24_U.if_read;
    assign fifo_intf_25.wr_en = AESL_inst_LINEAR.weights_stream_V_V_24_U.if_write;
    assign fifo_intf_25.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_024_blk_n);
    assign fifo_intf_25.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_094_blk_n);
    assign fifo_intf_25.finish = finish;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_LINEAR.weights_stream_V_V_25_U.if_read;
    assign fifo_intf_26.wr_en = AESL_inst_LINEAR.weights_stream_V_V_25_U.if_write;
    assign fifo_intf_26.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_025_blk_n);
    assign fifo_intf_26.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_095_blk_n);
    assign fifo_intf_26.finish = finish;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_LINEAR.weights_stream_V_V_26_U.if_read;
    assign fifo_intf_27.wr_en = AESL_inst_LINEAR.weights_stream_V_V_26_U.if_write;
    assign fifo_intf_27.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_026_blk_n);
    assign fifo_intf_27.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_096_blk_n);
    assign fifo_intf_27.finish = finish;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_LINEAR.weights_stream_V_V_27_U.if_read;
    assign fifo_intf_28.wr_en = AESL_inst_LINEAR.weights_stream_V_V_27_U.if_write;
    assign fifo_intf_28.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_027_blk_n);
    assign fifo_intf_28.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_097_blk_n);
    assign fifo_intf_28.finish = finish;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_LINEAR.weights_stream_V_V_28_U.if_read;
    assign fifo_intf_29.wr_en = AESL_inst_LINEAR.weights_stream_V_V_28_U.if_write;
    assign fifo_intf_29.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_028_blk_n);
    assign fifo_intf_29.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_098_blk_n);
    assign fifo_intf_29.finish = finish;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_LINEAR.weights_stream_V_V_29_U.if_read;
    assign fifo_intf_30.wr_en = AESL_inst_LINEAR.weights_stream_V_V_29_U.if_write;
    assign fifo_intf_30.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_029_blk_n);
    assign fifo_intf_30.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_099_blk_n);
    assign fifo_intf_30.finish = finish;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_LINEAR.weights_stream_V_V_30_U.if_read;
    assign fifo_intf_31.wr_en = AESL_inst_LINEAR.weights_stream_V_V_30_U.if_write;
    assign fifo_intf_31.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_030_blk_n);
    assign fifo_intf_31.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0100_blk_n);
    assign fifo_intf_31.finish = finish;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_LINEAR.weights_stream_V_V_31_U.if_read;
    assign fifo_intf_32.wr_en = AESL_inst_LINEAR.weights_stream_V_V_31_U.if_write;
    assign fifo_intf_32.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_031_blk_n);
    assign fifo_intf_32.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0101_blk_n);
    assign fifo_intf_32.finish = finish;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_LINEAR.iacts_stream_U.if_read;
    assign fifo_intf_33.wr_en = AESL_inst_LINEAR.iacts_stream_U.if_write;
    assign fifo_intf_33.fifo_rd_block = ~(AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.iacts_stream_blk_n);
    assign fifo_intf_33.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.iacts_stream64_blk_n);
    assign fifo_intf_33.finish = finish;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_LINEAR.X_c_U.if_read;
    assign fifo_intf_34.wr_en = AESL_inst_LINEAR.X_c_U.if_write;
    assign fifo_intf_34.fifo_rd_block = ~(AESL_inst_LINEAR.OutputBuffer_U0.X_blk_n);
    assign fifo_intf_34.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.X_c_blk_n);
    assign fifo_intf_34.finish = finish;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_LINEAR.Wt_Y_c_U.if_read;
    assign fifo_intf_35.wr_en = AESL_inst_LINEAR.Wt_Y_c_U.if_write;
    assign fifo_intf_35.fifo_rd_block = ~(AESL_inst_LINEAR.OutputBuffer_U0.Wt_Y_blk_n);
    assign fifo_intf_35.fifo_wr_block = ~(AESL_inst_LINEAR.ReadFromMem_U0.Wt_Y_c_blk_n);
    assign fifo_intf_35.finish = finish;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_LINEAR.block_num_x_loc_channel_U.if_read;
    assign fifo_intf_36.wr_en = AESL_inst_LINEAR.block_num_x_loc_channel_U.if_write;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_LINEAR.block_num_y_cast_loc_channel_U.if_read;
    assign fifo_intf_37.wr_en = AESL_inst_LINEAR.block_num_y_cast_loc_channel_U.if_write;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_LINEAR.ifc7_c_channel_U.if_read;
    assign fifo_intf_38.wr_en = AESL_inst_LINEAR.ifc7_c_channel_U.if_write;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;

    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_LINEAR.entry_proc_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_LINEAR.entry_proc_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_LINEAR.entry_proc_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_LINEAR.entry_proc_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_LINEAR.entry_proc_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.finish = finish;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_LINEAR.Block_split10_proc_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_LINEAR.Block_split10_proc_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_LINEAR.Block_split10_proc_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_LINEAR.Block_split10_proc_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_LINEAR.Block_split10_proc_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0;
    assign process_intf_2.finish = finish;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_LINEAR.ReadFromMem_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_LINEAR.ReadFromMem_U0.ap_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_071_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_072_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_073_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_074_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_075_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_076_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_077_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_078_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_079_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_080_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_081_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_082_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_083_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_084_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_085_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_086_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_087_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_088_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_089_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_090_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_091_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_092_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_093_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_094_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_095_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_096_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_097_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_098_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_099_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0100_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.weights_stream_0_0_0_0101_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.iacts_stream64_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.X_c_blk_n | ~AESL_inst_LINEAR.ReadFromMem_U0.Wt_Y_c_blk_n;
    assign process_intf_3.finish = finish;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_LINEAR.RunDataFlow_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_LINEAR.RunDataFlow_U0.ap_start;
    assign process_intf_4.pin_stall = 1'b0 | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.iacts_stream_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_0_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_01_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_02_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_03_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_04_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_05_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_06_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_07_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_08_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_09_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_010_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_011_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_012_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_013_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_014_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_015_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_016_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_017_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_018_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_019_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_020_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_021_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_022_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_023_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_024_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_025_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_026_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_027_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_028_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_029_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_030_blk_n | ~AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.weights_stream_0_0_0_031_blk_n;
    assign process_intf_4.pout_stall = 1'b0;
    assign process_intf_4.finish = finish;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_LINEAR.OutputBuffer_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_LINEAR.OutputBuffer_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_LINEAR.OutputBuffer_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_LINEAR.OutputBuffer_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_LINEAR.OutputBuffer_U0.ap_start;
    assign process_intf_5.pin_stall = 1'b0 | ~AESL_inst_LINEAR.OutputBuffer_U0.X_blk_n | ~AESL_inst_LINEAR.OutputBuffer_U0.Wt_Y_blk_n;
    assign process_intf_5.pout_stall = 1'b0;
    assign process_intf_5.finish = finish;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_LINEAR.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_LINEAR.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_LINEAR.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_230_2_fu_114.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_230_2_fu_114.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_230_2_fu_114.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_287_1_fu_67.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_287_1_fu_67.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_287_1_fu_67.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.grp_DPEUnit_fu_63.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.grp_DPEUnit_fu_63.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.grp_DPEUnit_fu_63.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;

    seq_loop_intf#(29) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b1;
    assign seq_loop_intf_1.one_state_block = AESL_inst_LINEAR.ReadFromMem_U0.ap_ST_fsm_state6_blk;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(29) seq_loop_monitor_1;
    seq_loop_intf#(6) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(6) seq_loop_monitor_2;
    seq_loop_intf#(6) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_LINEAR.RunDataFlow_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(6) seq_loop_monitor_3;
    seq_loop_intf#(4) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ST_fsm_state1;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ST_fsm_state4;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ST_fsm_state2;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ST_fsm_state2;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.ap_ST_fsm_state3;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(4) seq_loop_monitor_4;
    upc_loop_intf#(4) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_1.quit_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_1.loop_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_27_1_VITIS_LOOP_32_2_fu_576.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(4) upc_loop_monitor_1;
    upc_loop_intf#(12) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_ST_fsm_pp0_stage8;
    assign upc_loop_intf_2.quit_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_ST_fsm_pp0_stage8;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_block_pp0_stage8_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_block_pp0_stage8_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.loop_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_153_8_fu_747.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(12) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.loop_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_168_11_VITIS_LOOP_177_13_fu_757.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(20) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_ST_fsm_pp0_stage19;
    assign upc_loop_intf_4.quit_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_ST_fsm_pp0_stage19;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_block_pp0_stage19_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_block_pp0_stage19_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.quit_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_187_14_VITIS_LOOP_189_15_VITIS_LOOP_192_16_fu_767.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(20) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.loop_start = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_LINEAR.ReadFromMem_U0.grp_ReadFromMem_Pipeline_VITIS_LOOP_216_18_fu_980.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b0;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_CreateBitMask_fu_171.grp_CreateBitMask_Pipeline_VITIS_LOOP_237_3_VITIS_LOOP_241_4_fu_183.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.loop_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_RunDataFlow_Pipeline_VITIS_LOOP_341_1_fu_243.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b0;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.loop_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_291_2_fu_58.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b0;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(40) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.loop_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_296_3_fu_73.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b0;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(40) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.loop_start = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_LINEAR.RunDataFlow_U0.grp_DPEComputation_fu_250.grp_DPEComputation_Pipeline_VITIS_LOOP_303_4_fu_84.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b0;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(2) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_11.quit_state = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_LINEAR.OutputBuffer_U0.grp_OutputBuffer_Pipeline_VITIS_LOOP_329_1_fu_85.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b0;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(2) upc_loop_monitor_11;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
